sekundy_inst : sekundy PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
